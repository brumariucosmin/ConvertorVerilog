`ifndef __spi_intf
`define __spi_intf

interface spi_interface_dut;
  logic        sclk;
  logic        mosi;
  logic        miso;
  logic        cs;

 import uvm_pkg::*;
      
//ASERTII
      
endinterface


`endif