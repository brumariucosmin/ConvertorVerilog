`ifndef __button_intf
`define __button_intf

interface button_interface_dut;
  logic clk_i; 
  logic reset_n;
  logic enable_i;

endinterface

`endif