module apb_slave(pclk_i, rst_n_i, psel_i, penable_i, paddr_i);

  input pclk_i;
  input rst_n_i;
  input [2:0] paddr_i;
  input psel_i;
  input penable_i;

endmodule